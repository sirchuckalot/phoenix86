module (
  // We can optionally declare parameters here
  parameter <parameter_name> = <default_value>
)
cpu_top (
  // All IO are defined here
  <direction> <data_type> <size> <port_name>
);
 // Functional RTL (or structural) code
endmodule
